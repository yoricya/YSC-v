module ysc_interpreter

